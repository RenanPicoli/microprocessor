--------------------------------------------------
--instruction memory implementation
--by Renan Picoli de Souza
--supports only 32 bit instructions
--(all instructions are word-aligned)
--1024 bytes de ROM (como um I-cache)
--------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;--to_integer

use std.textio.all;--for file reading
use ieee.std_logic_textio.all;--for reading of std_logic_vectors

use work.my_types.all;--opcode and register "defines"

entity mini_rom is
	port (CLK: in std_logic;--borda de subida para escrita, se desativado, memória é lida
			RST: in std_logic;--asynchronous reset
			--interface de instrução (read-only)
			ADDR_A: in std_logic_vector(9 downto 0);--addr é endereço de byte, mas os Lsb são 00
			Q_A:	out std_logic_vector(31 downto 0);
			--interface de dados (read-write)
			D_B:	in std_logic_vector(31 downto 0);
			ADDR_B: in std_logic_vector(9 downto 0);--addr é endereço de byte, mas os Lsb são 00
			WREN_B: std_logic;
			Q_B:	out std_logic_vector(31 downto 0)
			);
end mini_rom;

architecture memArch of mini_rom is

	signal ADDR_reg_A: std_logic_vector((ADDR_A'length)-1 downto 0);--ADDR_A is registered, then it is used to select instruction
	signal ADDR_reg_B: std_logic_vector((ADDR_B'length)-1 downto 0);--ADDR_B is registered, then it is used to select instruction

	type memory is array (0 to 2**(ADDR_A'length)-1) of std_logic_vector(31 downto 0);
	constant initial_value: memory := (
0=> x"00000027",
1=> x"CFE00000",
2=> x"C3C00000",
3=> x"D400002E",
4=> x"C4400000",
5=> x"C8000000",
6=> x"D400004F",
7=> x"C4400000",
8=> x"C8000000",
9=> x"20040000",
10=> x"CC800000",
11=> x"D4000252",
12=> x"C4400000",
13=> x"C8000001",
14=> x"44400000",
15=> x"04420004",
16=> x"AFC2FFFB",
17=> x"44400000",
18=> x"04420030",
19=> x"AFC2FFFC",
20=> x"AFC0FFFD",
21=> x"23C2001C",
22=> x"20440000",
23=> x"CC800000",
24=> x"D40002A3",
25=> x"C4400000",
26=> x"C8000001",
27=> x"44800000",
28=> x"0484006A",
29=> x"CC800000",
30=> x"D400014B",
31=> x"C4400000",
32=> x"C8000001",
33=> x"AFC2FFFA",
34=> x"CC800000",
35=> x"D4000064",
36=> x"C4400000",
37=> x"C8000001",
38=> x"44800000",
39=> x"04840001",
40=> x"CC800000",
41=> x"D4000252",
42=> x"C4400000",
43=> x"C8000001",
44=> x"18000000",
45=> x"0800002C",
46=> x"00000027",
47=> x"00210827",
48=> x"00421027",
49=> x"00631827",
50=> x"00842027",
51=> x"00A52827",
52=> x"00C63027",
53=> x"00E73827",
54=> x"01084027",
55=> x"01294827",
56=> x"014A5027",
57=> x"016B5827",
58=> x"018C6027",
59=> x"01AD6827",
60=> x"01CE7027",
61=> x"01EF7827",
62=> x"02108027",
63=> x"02318827",
64=> x"02529027",
65=> x"02739827",
66=> x"0294A027",
67=> x"02B5A827",
68=> x"02D6B027",
69=> x"02F7B827",
70=> x"0318C027",
71=> x"0339C827",
72=> x"035AD027",
73=> x"037BD827",
74=> x"039CE027",
75=> x"03BDE827",
76=> x"03DEF027",
77=> x"03FFF827",
78=> x"D8000000",
79=> x"C3C00000",
80=> x"44400000",
81=> x"044200D0",
82=> x"AC0200A0",
83=> x"20020000",
84=> x"AC0200C0",
85=> x"44400000",
86=> x"04420100",
87=> x"AC0200A3",
88=> x"44400000",
89=> x"04420003",
90=> x"AC0200C1",
91=> x"44400000",
92=> x"044200F9",
93=> x"AC0200A1",
94=> x"44400000",
95=> x"04420001",
96=> x"AC0200C2",
97=> x"FC000000",
98=> x"CC400000",
99=> x"D8000000",
100=> x"CFE00000",
101=> x"C3C00000",
102=> x"44400000",
103=> x"04420100",
104=> x"AFC2FFFC",
105=> x"44400000",
106=> x"04420001",
107=> x"AFC2FFFD",
108=> x"23C20018",
109=> x"20440000",
110=> x"CC800000",
111=> x"D4000262",
112=> x"C4400000",
113=> x"C8000001",
114=> x"44A00000",
115=> x"04A51E00",
116=> x"44800000",
117=> x"0484001A",
118=> x"CCA00000",
119=> x"CC800000",
120=> x"D4000278",
121=> x"C4400000",
122=> x"C8000002",
123=> x"44A00000",
124=> x"04A50C77",
125=> x"44800000",
126=> x"0484001A",
127=> x"CCA00000",
128=> x"CC800000",
129=> x"D4000278",
130=> x"C4400000",
131=> x"C8000002",
132=> x"44A00000",
133=> x"04A50812",
134=> x"44800000",
135=> x"0484001A",
136=> x"CCA00000",
137=> x"CC800000",
138=> x"D4000278",
139=> x"C4400000",
140=> x"C8000002",
141=> x"44A00000",
142=> x"04A50A00",
143=> x"44800000",
144=> x"0484001A",
145=> x"CCA00000",
146=> x"CC800000",
147=> x"D4000278",
148=> x"C4400000",
149=> x"C8000002",
150=> x"44A00000",
151=> x"04A50E12",
152=> x"44800000",
153=> x"0484001A",
154=> x"CCA00000",
155=> x"CC800000",
156=> x"D4000278",
157=> x"C4400000",
158=> x"C8000002",
159=> x"44A00000",
160=> x"04A51023",
161=> x"44800000",
162=> x"0484001A",
163=> x"CCA00000",
164=> x"CC800000",
165=> x"D4000278",
166=> x"C4400000",
167=> x"C8000002",
168=> x"44A00000",
169=> x"04A50451",
170=> x"44800000",
171=> x"0484001A",
172=> x"CCA00000",
173=> x"CC800000",
174=> x"D4000278",
175=> x"C4400000",
176=> x"C8000002",
177=> x"44A00000",
178=> x"04A50651",
179=> x"44800000",
180=> x"0484001A",
181=> x"CCA00000",
182=> x"CC800000",
183=> x"D4000278",
184=> x"C4400000",
185=> x"C8000002",
186=> x"44A00000",
187=> x"04A51201",
188=> x"44800000",
189=> x"0484001A",
190=> x"CCA00000",
191=> x"CC800000",
192=> x"D4000278",
193=> x"C4400000",
194=> x"C8000002",
195=> x"44A00000",
196=> x"04A50C67",
197=> x"44800000",
198=> x"0484001A",
199=> x"CCA00000",
200=> x"CC800000",
201=> x"D4000278",
202=> x"C4400000",
203=> x"C8000002",
204=> x"FC000000",
205=> x"D3E00000",
206=> x"CC400000",
207=> x"D8000000",
208=> x"CFE00000",
209=> x"C3C00000",
210=> x"1C000258",
211=> x"8C020030",
212=> x"AFC2FFFB",
213=> x"8FC2FFFB",
214=> x"20450000",
215=> x"44800000",
216=> x"8C840705",
217=> x"CCA00000",
218=> x"CC800000",
219=> x"D40002F9",
220=> x"C4400000",
221=> x"C8000002",
222=> x"20430000",
223=> x"44400000",
224=> x"8C420706",
225=> x"20450000",
226=> x"20640000",
227=> x"CCA00000",
228=> x"CC800000",
229=> x"D4000126",
230=> x"C4400000",
231=> x"C8000002",
232=> x"AFC2FFFA",
233=> x"44400000",
234=> x"8C420707",
235=> x"8FC3FFFA",
236=> x"00421801",
237=> x"AFC2FFFC",
238=> x"8FC2FFFC",
239=> x"AC020010",
240=> x"8C020071",
241=> x"AFC2FFFD",
242=> x"8FC2FFFD",
243=> x"AC020011",
244=> x"DC000000",
245=> x"FC000000",
246=> x"D3E00000",
247=> x"CC400000",
248=> x"D8000000",
249=> x"C3C00000",
250=> x"20020000",
251=> x"AC020064",
252=> x"DC000000",
253=> x"FC000000",
254=> x"CC400000",
255=> x"D8000000",
256=> x"C3C00000",
257=> x"8C020070",
258=> x"AFC2FFF8",
259=> x"8C020011",
260=> x"AFC2FFF9",
261=> x"8FC2FFF9",
262=> x"8FC3FFF8",
263=> x"00421802",
264=> x"AFC2FFFA",
265=> x"8C020010",
266=> x"AFC2FFFB",
267=> x"8FC2FFFB",
268=> x"8FC3FFFA",
269=> x"00421801",
270=> x"AFC2FFFC",
271=> x"8FC2FFFC",
272=> x"AC020050",
273=> x"1C000020",
274=> x"3C000000",
275=> x"1C000501",
276=> x"1C000002",
277=> x"8C020073",
278=> x"AFC2FFF6",
279=> x"8FC2FFF6",
280=> x"AC020069",
281=> x"8FC2FFF6",
282=> x"AC020069",
283=> x"8C020068",
284=> x"AFC2FFF7",
285=> x"8FC2FFF7",
286=> x"04420001",
287=> x"AFC2FFF7",
288=> x"8FC2FFF7",
289=> x"AC020068",
290=> x"DC000000",
291=> x"FC000000",
292=> x"CC400000",
293=> x"D8000000",
294=> x"CFE00000",
295=> x"C3C00000",
296=> x"8FC50001",
297=> x"8FC40000",
298=> x"CCA00000",
299=> x"CC800000",
300=> x"D40002ED",
301=> x"C4400000",
302=> x"C8000002",
303=> x"AFC2FFFC",
304=> x"8FC3FFFC",
305=> x"44408000",
306=> x"04420000",
307=> x"00621024",
308=> x"AFC2FFFC",
309=> x"8FC3FFFC",
310=> x"44408000",
311=> x"04420000",
312=> x"10620001",
313=> x"0800013C",
314=> x"8FC20000",
315=> x"0800013D",
316=> x"8FC20001",
317=> x"D3E00000",
318=> x"CC400000",
319=> x"D8000000",
320=> x"C0400000",
321=> x"8C410000",
322=> x"00631827",
323=> x"20630074",
324=> x"AC610000",
325=> x"D8000000",
326=> x"C0400000",
327=> x"8C410001",
328=> x"8C440000",
329=> x"AC810000",
330=> x"D8000000",
331=> x"C3C00000",
332=> x"8FC40000",
333=> x"8C820000",
334=> x"CC400000",
335=> x"D8000000",
336=> x"C3C00000",
337=> x"8FC40000",
338=> x"8FC50001",
339=> x"8FC60002",
340=> x"00210827",
341=> x"00811020",
342=> x"00A11820",
343=> x"8C480000",
344=> x"AC680000",
345=> x"20210001",
346=> x"10260001",
347=> x"08000155",
348=> x"D8000000",
349=> x"C3C00000",
350=> x"8FC40000",
351=> x"8FC50001",
352=> x"00C63027",
353=> x"20C60008",
354=> x"00210827",
355=> x"00811020",
356=> x"00A11820",
357=> x"8C480000",
358=> x"AC680000",
359=> x"20210001",
360=> x"10260001",
361=> x"08000155",
362=> x"D8000000",
363=> x"CFE00000",
364=> x"C3C00000",
365=> x"8FC60002",
366=> x"44A00000",
367=> x"04A50020",
368=> x"8FC40000",
369=> x"CCC00000",
370=> x"CCA00000",
371=> x"CC800000",
372=> x"D4000150",
373=> x"C4400000",
374=> x"C8000003",
375=> x"8FC60002",
376=> x"44A00000",
377=> x"04A50028",
378=> x"8FC40001",
379=> x"CCC00000",
380=> x"CCA00000",
381=> x"CC800000",
382=> x"D4000150",
383=> x"C4400000",
384=> x"C8000003",
385=> x"44800000",
386=> x"04840030",
387=> x"CCC00000",
388=> x"CCA00000",
389=> x"CC800000",
390=> x"D400014B",
391=> x"C4400000",
392=> x"C8000003",
393=> x"AFC2FFFC",
394=> x"8FC2FFFC",
395=> x"D3E00000",
396=> x"CC400000",
397=> x"D8000000",
398=> x"CFE00000",
399=> x"C3C00000",
400=> x"44A00000",
401=> x"04A50040",
402=> x"8FC40000",
403=> x"CCC00000",
404=> x"CCA00000",
405=> x"CC800000",
406=> x"D400015D",
407=> x"C4400000",
408=> x"C8000003",
409=> x"44A00000",
410=> x"04A50048",
411=> x"8FC40001",
412=> x"CCC00000",
413=> x"CCA00000",
414=> x"CC800000",
415=> x"D400015D",
416=> x"C4400000",
417=> x"C8000003",
418=> x"8FC50002",
419=> x"44800000",
420=> x"04840050",
421=> x"CCC00000",
422=> x"CCA00000",
423=> x"CC800000",
424=> x"D4000146",
425=> x"C4400000",
426=> x"C8000003",
427=> x"3C000000",
428=> x"8FC50000",
429=> x"44800000",
430=> x"04840040",
431=> x"CCC00000",
432=> x"CCA00000",
433=> x"CC800000",
434=> x"D400015D",
435=> x"C4400000",
436=> x"C8000003",
437=> x"FC000000",
438=> x"D3E00000",
439=> x"CC400000",
440=> x"D8000000",
441=> x"CFE00000",
442=> x"CE000000",
443=> x"C3C00000",
444=> x"AFC70003",
445=> x"AFC0FFFA",
446=> x"080001DE",
447=> x"8FC30004",
448=> x"8FC2FFFA",
449=> x"00628020",
450=> x"8FC3FFFA",
451=> x"8FC20003",
452=> x"34620000",
453=> x"94600000",
454=> x"8FC20000",
455=> x"00621020",
456=> x"8FC60003",
457=> x"8FC50002",
458=> x"20440000",
459=> x"CCE00000",
460=> x"CCC00000",
461=> x"CCA00000",
462=> x"CC800000",
463=> x"D400016B",
464=> x"C4400000",
465=> x"C8000004",
466=> x"20450000",
467=> x"22040000",
468=> x"CCE00000",
469=> x"CCC00000",
470=> x"CCA00000",
471=> x"CC800000",
472=> x"D4000146",
473=> x"C4400000",
474=> x"C8000004",
475=> x"8FC2FFFA",
476=> x"20420001",
477=> x"AFC2FFFA",
478=> x"8FC3FFFA",
479=> x"8FC20001",
480=> x"00621022",
481=> x"004207D3",
482=> x"10400001",
483=> x"080001BF",
484=> x"FC000000",
485=> x"D3E00000",
486=> x"D2000000",
487=> x"CC400000",
488=> x"D8000000",
489=> x"CFE00000",
490=> x"C3C00000",
491=> x"AFC0FFF8",
492=> x"08000248",
493=> x"AFC0FFF9",
494=> x"0800023F",
495=> x"8FC60003",
496=> x"44A00000",
497=> x"04A50020",
498=> x"8FC40000",
499=> x"CCE00000",
500=> x"CCC00000",
501=> x"CCA00000",
502=> x"CC800000",
503=> x"D4000150",
504=> x"C4400000",
505=> x"C8000004",
506=> x"AFC0FFFA",
507=> x"0800021B",
508=> x"8FC30001",
509=> x"8FC2FFF9",
510=> x"00621820",
511=> x"8FC4FFFA",
512=> x"8FC20004",
513=> x"34820000",
514=> x"94400000",
515=> x"00621020",
516=> x"20440000",
517=> x"CCE00000",
518=> x"CCC00000",
519=> x"CCA00000",
520=> x"CC800000",
521=> x"D400014B",
522=> x"C4400000",
523=> x"C8000004",
524=> x"AFC2FFFC",
525=> x"8FC2FFFA",
526=> x"20420048",
527=> x"8FC5FFFC",
528=> x"20440000",
529=> x"CCE00000",
530=> x"CCC00000",
531=> x"CCA00000",
532=> x"CC800000",
533=> x"D4000146",
534=> x"C4400000",
535=> x"C8000004",
536=> x"8FC2FFFA",
537=> x"20420001",
538=> x"AFC2FFFA",
539=> x"8FC3FFFA",
540=> x"8FC20003",
541=> x"00621022",
542=> x"004207D3",
543=> x"10400001",
544=> x"080001FC",
545=> x"44800000",
546=> x"04840030",
547=> x"CCE00000",
548=> x"CCC00000",
549=> x"CCA00000",
550=> x"CC800000",
551=> x"D400014B",
552=> x"C4400000",
553=> x"C8000004",
554=> x"AFC2FFFB",
555=> x"8FC3FFF8",
556=> x"8FC20004",
557=> x"34620000",
558=> x"94600000",
559=> x"8FC20005",
560=> x"00621820",
561=> x"8FC2FFF9",
562=> x"00621020",
563=> x"8FC5FFFB",
564=> x"20440000",
565=> x"CCE00000",
566=> x"CCC00000",
567=> x"CCA00000",
568=> x"CC800000",
569=> x"D4000146",
570=> x"C4400000",
571=> x"C8000004",
572=> x"8FC2FFF9",
573=> x"20420001",
574=> x"AFC2FFF9",
575=> x"8FC3FFF9",
576=> x"8FC20004",
577=> x"00621022",
578=> x"004207D3",
579=> x"10400001",
580=> x"080001EF",
581=> x"8FC2FFF8",
582=> x"20420001",
583=> x"AFC2FFF8",
584=> x"8FC3FFF8",
585=> x"8FC20002",
586=> x"00621022",
587=> x"004207D3",
588=> x"10400001",
589=> x"080001ED",
590=> x"FC000000",
591=> x"D3E00000",
592=> x"CC400000",
593=> x"D8000000",
594=> x"CFE00000",
595=> x"C3C00000",
596=> x"8FC50000",
597=> x"44800000",
598=> x"04840072",
599=> x"CCE00000",
600=> x"CCC00000",
601=> x"CCA00000",
602=> x"CC800000",
603=> x"D4000146",
604=> x"C4400000",
605=> x"C8000004",
606=> x"FC000000",
607=> x"D3E00000",
608=> x"CC400000",
609=> x"D8000000",
610=> x"CFE00000",
611=> x"C3C00000",
612=> x"8FC20000",
613=> x"8C430000",
614=> x"8FC20000",
615=> x"8C420004",
616=> x"00621025",
617=> x"AFC2FFFC",
618=> x"8FC5FFFC",
619=> x"44800000",
620=> x"04840060",
621=> x"CCE00000",
622=> x"CCC00000",
623=> x"CCA00000",
624=> x"CC800000",
625=> x"D4000146",
626=> x"C4400000",
627=> x"C8000004",
628=> x"FC000000",
629=> x"D3E00000",
630=> x"CC400000",
631=> x"D8000000",
632=> x"CFE00000",
633=> x"C3C00000",
634=> x"8FC50001",
635=> x"44800000",
636=> x"04840061",
637=> x"CCE00000",
638=> x"CCC00000",
639=> x"CCA00000",
640=> x"CC800000",
641=> x"D4000146",
642=> x"C4400000",
643=> x"C8000004",
644=> x"44800000",
645=> x"04840060",
646=> x"CCE00000",
647=> x"CCC00000",
648=> x"CCA00000",
649=> x"CC800000",
650=> x"D400014B",
651=> x"C4400000",
652=> x"C8000004",
653=> x"AFC2FFFC",
654=> x"8FC20000",
655=> x"00430052",
656=> x"8FC2FFFC",
657=> x"00621025",
658=> x"04420400",
659=> x"AFC2FFFC",
660=> x"8FC5FFFC",
661=> x"44800000",
662=> x"04840060",
663=> x"CCE00000",
664=> x"CCC00000",
665=> x"CCA00000",
666=> x"CC800000",
667=> x"D4000146",
668=> x"C4400000",
669=> x"C8000004",
670=> x"18000000",
671=> x"FC000000",
672=> x"D3E00000",
673=> x"CC400000",
674=> x"D8000000",
675=> x"CFE00000",
676=> x"C3C00000",
677=> x"8FC20000",
678=> x"8C430008",
679=> x"8FC20000",
680=> x"8C420000",
681=> x"00621025",
682=> x"AFC2FFFC",
683=> x"8FC5FFFC",
684=> x"44800000",
685=> x"04840068",
686=> x"CCE00000",
687=> x"CCC00000",
688=> x"CCA00000",
689=> x"CC800000",
690=> x"D4000146",
691=> x"C4400000",
692=> x"C8000004",
693=> x"FC000000",
694=> x"D3E00000",
695=> x"CC400000",
696=> x"D8000000",
697=> x"CFE00000",
698=> x"C3C00000",
699=> x"8FC50001",
700=> x"44800000",
701=> x"04840069",
702=> x"CCE00000",
703=> x"CCC00000",
704=> x"CCA00000",
705=> x"CC800000",
706=> x"D4000146",
707=> x"C4400000",
708=> x"C8000004",
709=> x"44800000",
710=> x"04840068",
711=> x"CCE00000",
712=> x"CCC00000",
713=> x"CCA00000",
714=> x"CC800000",
715=> x"D400014B",
716=> x"C4400000",
717=> x"C8000004",
718=> x"AFC2FFFC",
719=> x"8FC2FFFC",
720=> x"04420003",
721=> x"AFC2FFFC",
722=> x"8FC5FFFC",
723=> x"44800000",
724=> x"04840068",
725=> x"CCE00000",
726=> x"CCC00000",
727=> x"CCA00000",
728=> x"CC800000",
729=> x"D4000146",
730=> x"C4400000",
731=> x"C8000004",
732=> x"FC000000",
733=> x"D3E00000",
734=> x"CC400000",
735=> x"D8000000",
736=> x"C3C00000",
737=> x"44600000",
738=> x"04630001",
739=> x"8FC20000",
740=> x"00621016",
741=> x"CC400000",
742=> x"D8000000",
743=> x"C0400000",
744=> x"8C430000",
745=> x"8C440001",
746=> x"00640800",
747=> x"CC200000",
748=> x"D8000000",
749=> x"C0400000",
750=> x"8C430000",
751=> x"8C440001",
752=> x"00640802",
753=> x"CC200000",
754=> x"D8000000",
755=> x"C0400000",
756=> x"8C430000",
757=> x"8C440001",
758=> x"00640801",
759=> x"CC200000",
760=> x"D8000000",
761=> x"C0400000",
762=> x"8C430000",
763=> x"8C440001",
764=> x"00640803",
765=> x"CC200000",
766=> x"D8000000",
767=> x"C0400000",
768=> x"8C430000",
769=> x"44808000",
770=> x"00641827",
771=> x"CC600000",
772=> x"D8000000",
773=> x"3F000000",
774=> x"461C4000",
775=> x"40000000",
others=> x"00000000"

	);
	signal rom: memory := initial_value;

	begin
		--output behaviour:
		--necessary turn Auto ROM Replacement on
		process(CLK,RST,ADDR_A)
		begin
--			if(RST='1')then
--				ADDR_reg_A <= (others=>'0');
			if(rising_edge(CLK))then
--				ADDR_reg_A <= ADDR_A;				
				Q_A <= rom(to_integer(unsigned(ADDR_A)));
			end if;
		end process;
		--surprisingly, the design also works with the synchronous reading logic (ram inferrence)
--		Q_A <= rom(to_integer(unsigned(ADDR_reg_A)));
--		Q_A <= rom(to_integer(unsigned(ADDR_A)));
		
		process(CLK,RST,ADDR_B,WREN_B)
		begin
--			if(RST='1')then
--				ADDR_reg_B <= (others=>'0');
--				rom <= initial_value;
--			elsif(rising_edge(CLK) and WREN_B='1')then
			if(rising_edge(CLK))then
--				ADDR_reg_B <= ADDR_B;
				if(WREN_B='1')then
					rom(to_integer(unsigned(ADDR_B))) <= D_B;
				end if;
				Q_B <= rom(to_integer(unsigned(ADDR_B)));
			end if;
		end process;		
		--surprisingly, the design also works with the synchronous reading logic (ram inferrence)
--		Q_B <= rom(to_integer(unsigned(ADDR_reg_B)));
--		Q_B <= rom(to_integer(unsigned(ADDR_B)));
end memArch;
