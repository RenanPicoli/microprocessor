--------------------------------------------------
--instruction memory implementation
--by Renan Picoli de Souza
--supports only 32 bit instructions
--(all instructions are word-aligned)
--1024 bytes de ROM (como um I-cache)
--------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;--to_integer

use std.textio.all;--for file reading
use ieee.std_logic_textio.all;--for reading of std_logic_vectors

use work.my_types.all;--opcode and register "defines"

entity mini_rom is
	port (
			RST: in std_logic;--asynchronous reset
			--interface de instrução (read-only)
			CLK_A:in std_logic;--borda de subida para escrita, se desativado, memória é lida
			ADDR_A: in std_logic_vector;--addr é endereço de byte, mas os Lsb são 00
			Q_A:	out std_logic_vector(31 downto 0);
			--interface de dados (read-write)
			CLK_B:in std_logic;--borda de subida para escrita, se desativado, memória é lida
			D_B:	in std_logic_vector(31 downto 0);
			ADDR_B: in std_logic_vector;--addr é endereço de byte, mas os Lsb são 00
			WREN_B: std_logic;
			Q_B:	out std_logic_vector(31 downto 0)
			);
end mini_rom;

architecture memArch of mini_rom is

	signal ADDR_reg_A: std_logic_vector((ADDR_A'length)-1 downto 0);--ADDR_A is registered, then it is used to select instruction
	signal ADDR_reg_B: std_logic_vector((ADDR_B'length)-1 downto 0);--ADDR_B is registered, then it is used to select instruction

	type memory is array (0 to 2**(ADDR_A'length)-1) of std_logic_vector(31 downto 0);
	constant initial_value: memory := (
0=> x"00000027",
1=> x"C800FFC0",
2=> x"CFE00000",
3=> x"C3C00000",
4=> x"44400000",
5=> x"8C423A34",
6=> x"AFC2FFDC",
7=> x"44400000",
8=> x"8C423A38",
9=> x"AFC2FFE0",
10=> x"44400000",
11=> x"8C423A3C",
12=> x"AFC2FFE4",
13=> x"D400004D",
14=> x"C4400000",
15=> x"C8000004",
16=> x"20040000",
17=> x"CC800000",
18=> x"D4000280",
19=> x"C4400000",
20=> x"C8000008",
21=> x"44400000",
22=> x"04420004",
23=> x"AFC2FFE8",
24=> x"44400000",
25=> x"04420030",
26=> x"AFC2FFEC",
27=> x"AFC0FFF0",
28=> x"23C2FFE8",
29=> x"20440000",
30=> x"CC800000",
31=> x"D40002CB",
32=> x"C4400000",
33=> x"C8000008",
34=> x"44800000",
35=> x"048401A8",
36=> x"CC800000",
37=> x"D400017C",
38=> x"C4400000",
39=> x"C8000008",
40=> x"AFC2FFD8",
41=> x"0C420080",
42=> x"10400001",
43=> x"10000001",
44=> x"08000022",
45=> x"D400006E",
46=> x"C4400000",
47=> x"C8000004",
48=> x"8FC4FFDC",
49=> x"CC800000",
50=> x"D4000546",
51=> x"C4400000",
52=> x"C800000C",
53=> x"44400000",
54=> x"0442022C",
55=> x"AC0201D4",
56=> x"8FC4FFE0",
57=> x"CC800000",
58=> x"D4000546",
59=> x"C4400000",
60=> x"C800000C",
61=> x"44400000",
62=> x"0442022C",
63=> x"AC0201D4",
64=> x"8FC4FFE4",
65=> x"CC800000",
66=> x"D4000546",
67=> x"C4400000",
68=> x"C800000C",
69=> x"44800000",
70=> x"04840001",
71=> x"CC800000",
72=> x"D4000280",
73=> x"C4400000",
74=> x"C8000008",
75=> x"18000000",
76=> x"0800004B",
77=> x"C800FFF8",
78=> x"C3C00000",
79=> x"44400000",
80=> x"04422368",
81=> x"2042E000",
82=> x"AC020280",
83=> x"20020000",
84=> x"AC020300",
85=> x"44400000",
86=> x"04422408",
87=> x"2042E000",
88=> x"AC02028C",
89=> x"44400000",
90=> x"04420003",
91=> x"AC020304",
92=> x"44400000",
93=> x"044223FC",
94=> x"2042E000",
95=> x"AC020284",
96=> x"44400000",
97=> x"04420001",
98=> x"AC020308",
99=> x"44400000",
100=> x"0442254C",
101=> x"2042E000",
102=> x"AC020290",
103=> x"44400000",
104=> x"04420004",
105=> x"AC02037C",
106=> x"FC000000",
107=> x"C8000008",
108=> x"CC400000",
109=> x"D8000000",
110=> x"C800FFD8",
111=> x"CFE00000",
112=> x"C3C00000",
113=> x"44400000",
114=> x"04420100",
115=> x"AFC2FFF0",
116=> x"AFC0FFF4",
117=> x"23C2FFF0",
118=> x"20440000",
119=> x"CC800000",
120=> x"D4000290",
121=> x"C4400000",
122=> x"C8000008",
123=> x"44A00000",
124=> x"04A51E00",
125=> x"44800000",
126=> x"0484001A",
127=> x"CCA00000",
128=> x"CC800000",
129=> x"D40002A6",
130=> x"C4400000",
131=> x"C800000C",
132=> x"44A00000",
133=> x"04A50C77",
134=> x"44800000",
135=> x"0484001A",
136=> x"CCA00000",
137=> x"CC800000",
138=> x"D40002A6",
139=> x"C4400000",
140=> x"C800000C",
141=> x"44A00000",
142=> x"04A50812",
143=> x"44800000",
144=> x"0484001A",
145=> x"CCA00000",
146=> x"CC800000",
147=> x"D40002A6",
148=> x"C4400000",
149=> x"C800000C",
150=> x"44A00000",
151=> x"04A50A00",
152=> x"44800000",
153=> x"0484001A",
154=> x"CCA00000",
155=> x"CC800000",
156=> x"D40002A6",
157=> x"C4400000",
158=> x"C800000C",
159=> x"44A00000",
160=> x"04A50E12",
161=> x"44800000",
162=> x"0484001A",
163=> x"CCA00000",
164=> x"CC800000",
165=> x"D40002A6",
166=> x"C4400000",
167=> x"C800000C",
168=> x"44A00000",
169=> x"04A51023",
170=> x"44800000",
171=> x"0484001A",
172=> x"CCA00000",
173=> x"CC800000",
174=> x"D40002A6",
175=> x"C4400000",
176=> x"C800000C",
177=> x"44A00000",
178=> x"04A50451",
179=> x"44800000",
180=> x"0484001A",
181=> x"CCA00000",
182=> x"CC800000",
183=> x"D40002A6",
184=> x"C4400000",
185=> x"C800000C",
186=> x"44A00000",
187=> x"04A50651",
188=> x"44800000",
189=> x"0484001A",
190=> x"CCA00000",
191=> x"CC800000",
192=> x"D40002A6",
193=> x"C4400000",
194=> x"C800000C",
195=> x"44A00000",
196=> x"04A51201",
197=> x"44800000",
198=> x"0484001A",
199=> x"CCA00000",
200=> x"CC800000",
201=> x"D40002A6",
202=> x"C4400000",
203=> x"C800000C",
204=> x"44A00000",
205=> x"04A50C67",
206=> x"44800000",
207=> x"0484001A",
208=> x"CCA00000",
209=> x"CC800000",
210=> x"D40002A6",
211=> x"C4400000",
212=> x"C800000C",
213=> x"FC000000",
214=> x"D3E00000",
215=> x"C8000028",
216=> x"CC400000",
217=> x"D8000000",
218=> x"44400000",
219=> x"04420002",
220=> x"44600000",
221=> x"04630058",
222=> x"48430000",
223=> x"44400000",
224=> x"04420001",
225=> x"AC0200C4",
226=> x"8C0200C0",
227=> x"AFC2FFE4",
228=> x"20430000",
229=> x"44400000",
230=> x"8C423A40",
231=> x"00431003",
232=> x"AFC2FFE8",
233=> x"44400000",
234=> x"8C423A44",
235=> x"20450000",
236=> x"8FC4FFE8",
237=> x"CCA00000",
238=> x"CC800000",
239=> x"D4000154",
240=> x"C4400000",
241=> x"C800000C",
242=> x"AFC2FFE0",
243=> x"44400000",
244=> x"8C423A48",
245=> x"8FC3FFE0",
246=> x"00431001",
247=> x"AFC2FFEC",
248=> x"AC020040",
249=> x"8C0201C4",
250=> x"AFC2FFF0",
251=> x"AC020044",
252=> x"8FC2FFE4",
253=> x"AC020048",
254=> x"DC000000",
255=> x"20020000",
256=> x"AC020190",
257=> x"DC000000",
258=> x"8C0201C0",
259=> x"AFC2FFD0",
260=> x"8C020044",
261=> x"AFC2FFD4",
262=> x"8FC3FFD0",
263=> x"00431002",
264=> x"AFC2FFD8",
265=> x"8C020040",
266=> x"AFC2FFDC",
267=> x"8FC3FFD8",
268=> x"00431001",
269=> x"AFC2FFE0",
270=> x"AC020140",
271=> x"20030000",
272=> x"44400000",
273=> x"04420020",
274=> x"48620000",
275=> x"3C000000",
276=> x"44400000",
277=> x"04420005",
278=> x"44600000",
279=> x"04630001",
280=> x"48430000",
281=> x"20030000",
282=> x"44400000",
283=> x"0442001A",
284=> x"48620000",
285=> x"44400000",
286=> x"04420001",
287=> x"AC0200C4",
288=> x"8C0200C0",
289=> x"AFC2FFE4",
290=> x"8C0201CC",
291=> x"20500000",
292=> x"AC0201A4",
293=> x"AC0201A4",
294=> x"8C0201A0",
295=> x"20500000",
296=> x"04500001",
297=> x"AC1001A0",
298=> x"8FC2FFE0",
299=> x"8FC3FFE0",
300=> x"00431001",
301=> x"AFC2FFE8",
302=> x"8C020048",
303=> x"AFC2FFEC",
304=> x"8FC2FFE8",
305=> x"8FC3FFEC",
306=> x"00431001",
307=> x"AFC2FFEC",
308=> x"8FC3FFE4",
309=> x"00431003",
310=> x"20500000",
311=> x"44400000",
312=> x"8C423A4C",
313=> x"02021002",
314=> x"AFC2FFF0",
315=> x"CE000000",
316=> x"0040802A",
317=> x"12000002",
318=> x"D2000000",
319=> x"10000002",
320=> x"D2000000",
321=> x"08000152",
322=> x"44400000",
323=> x"8C423A54",
324=> x"10400001",
325=> x"08000152",
326=> x"44400000",
327=> x"04420001",
328=> x"44000000",
329=> x"AC023A54",
330=> x"00000027",
331=> x"20030000",
332=> x"44400000",
333=> x"04420080",
334=> x"48620000",
335=> x"44400000",
336=> x"04420010",
337=> x"AC020214",
338=> x"DC000000",
339=> x"DC000000",
340=> x"C800FFD8",
341=> x"CFE00000",
342=> x"C3C00000",
343=> x"AFC40000",
344=> x"AFC50004",
345=> x"8FC40000",
346=> x"CCA00000",
347=> x"CC800000",
348=> x"D4000314",
349=> x"C4400000",
350=> x"C800000C",
351=> x"AFC2FFF0",
352=> x"20430000",
353=> x"44408000",
354=> x"04420000",
355=> x"00621024",
356=> x"AFC2FFF0",
357=> x"20430000",
358=> x"44408000",
359=> x"04420000",
360=> x"10620001",
361=> x"0800016C",
362=> x"8FC20000",
363=> x"0800016D",
364=> x"8FC20004",
365=> x"D3E00000",
366=> x"C8000028",
367=> x"CC400000",
368=> x"D8000000",
369=> x"C0400000",
370=> x"8C410000",
371=> x"00631827",
372=> x"206301D0",
373=> x"AC610000",
374=> x"D8000000",
375=> x"C0400000",
376=> x"8C410004",
377=> x"8C440000",
378=> x"AC810000",
379=> x"D8000000",
380=> x"C3C00000",
381=> x"8FC40000",
382=> x"8C820000",
383=> x"CC400000",
384=> x"D8000000",
385=> x"C3C00000",
386=> x"8FC40000",
387=> x"8FC50004",
388=> x"8FC60008",
389=> x"00210827",
390=> x"00811020",
391=> x"00A11820",
392=> x"8C480000",
393=> x"AC680000",
394=> x"20210001",
395=> x"10260001",
396=> x"08000186",
397=> x"D8000000",
398=> x"C3C00000",
399=> x"8FC40000",
400=> x"8FC50004",
401=> x"00C63027",
402=> x"20C60008",
403=> x"00210827",
404=> x"00811020",
405=> x"00A11820",
406=> x"8C480000",
407=> x"AC680000",
408=> x"20210001",
409=> x"10260001",
410=> x"08000186",
411=> x"D8000000",
412=> x"C800FFD8",
413=> x"CFE00000",
414=> x"C3C00000",
415=> x"AFC40000",
416=> x"AFC50004",
417=> x"AFC60008",
418=> x"44A00000",
419=> x"04A50080",
420=> x"8FC40000",
421=> x"CCC00000",
422=> x"CCA00000",
423=> x"CC800000",
424=> x"D4000181",
425=> x"C800000C",
426=> x"8FC60008",
427=> x"44A00000",
428=> x"04A500A0",
429=> x"8FC40004",
430=> x"CCC00000",
431=> x"CCA00000",
432=> x"CC800000",
433=> x"D4000181",
434=> x"C800000C",
435=> x"44A00000",
436=> x"04A50001",
437=> x"44800000",
438=> x"048400C4",
439=> x"CCA00000",
440=> x"CC800000",
441=> x"D4000177",
442=> x"C8000008",
443=> x"44800000",
444=> x"048400C0",
445=> x"CC800000",
446=> x"D400017C",
447=> x"C4400000",
448=> x"C8000008",
449=> x"AFC2FFF0",
450=> x"D3E00000",
451=> x"C8000028",
452=> x"CC400000",
453=> x"D8000000",
454=> x"C800FFE0",
455=> x"CFE00000",
456=> x"C3C00000",
457=> x"AFC40000",
458=> x"AFC50004",
459=> x"AFC60008",
460=> x"44A00000",
461=> x"04A50100",
462=> x"8FC40000",
463=> x"CCA00000",
464=> x"CC800000",
465=> x"D400018E",
466=> x"C8000008",
467=> x"44A00000",
468=> x"04A50120",
469=> x"8FC40004",
470=> x"CCA00000",
471=> x"CC800000",
472=> x"D400018E",
473=> x"C8000008",
474=> x"8FC50008",
475=> x"44800000",
476=> x"04840140",
477=> x"CCA00000",
478=> x"CC800000",
479=> x"D4000177",
480=> x"C8000008",
481=> x"3C000000",
482=> x"8FC50000",
483=> x"44800000",
484=> x"04840100",
485=> x"CCA00000",
486=> x"CC800000",
487=> x"D400018E",
488=> x"C8000008",
489=> x"FC000000",
490=> x"D3E00000",
491=> x"C8000020",
492=> x"CC400000",
493=> x"D8000000",
494=> x"C800FFD0",
495=> x"CFE00000",
496=> x"CE000000",
497=> x"C3C00000",
498=> x"AFC40000",
499=> x"AFC50004",
500=> x"AFC60008",
501=> x"AFC7000C",
502=> x"AFC0FFE8",
503=> x"08000213",
504=> x"8FC30010",
505=> x"8FC2FFE8",
506=> x"00628020",
507=> x"8FC3FFE8",
508=> x"8FC2000C",
509=> x"34620000",
510=> x"94600000",
511=> x"8FC20000",
512=> x"00621020",
513=> x"8FC6000C",
514=> x"8FC50008",
515=> x"20440000",
516=> x"CCC00000",
517=> x"CCA00000",
518=> x"CC800000",
519=> x"D400019C",
520=> x"C4400000",
521=> x"C8000010",
522=> x"20450000",
523=> x"22040000",
524=> x"CCA00000",
525=> x"CC800000",
526=> x"D4000177",
527=> x"C8000008",
528=> x"8FC2FFE8",
529=> x"20420001",
530=> x"AFC2FFE8",
531=> x"8FC3FFE8",
532=> x"8FC20004",
533=> x"00621022",
534=> x"004207D3",
535=> x"10400001",
536=> x"080001F8",
537=> x"FC000000",
538=> x"D3E00000",
539=> x"D2000000",
540=> x"C8000030",
541=> x"CC400000",
542=> x"D8000000",
543=> x"C800FFC8",
544=> x"CFE00000",
545=> x"C3C00000",
546=> x"AFC40000",
547=> x"AFC50004",
548=> x"AFC60008",
549=> x"AFC7000C",
550=> x"AFC0FFE0",
551=> x"08000275",
552=> x"AFC0FFE4",
553=> x"0800026C",
554=> x"8FC6000C",
555=> x"44A00000",
556=> x"04A50080",
557=> x"8FC40000",
558=> x"CCC00000",
559=> x"CCA00000",
560=> x"CC800000",
561=> x"D4000181",
562=> x"C800000C",
563=> x"AFC0FFE8",
564=> x"0800024E",
565=> x"8FC30004",
566=> x"8FC2FFE4",
567=> x"00621820",
568=> x"8FC4FFE8",
569=> x"8FC20010",
570=> x"34820000",
571=> x"94400000",
572=> x"00621020",
573=> x"20440000",
574=> x"CC800000",
575=> x"D400017C",
576=> x"C4400000",
577=> x"C8000008",
578=> x"AFC2FFF0",
579=> x"8FC2FFE8",
580=> x"20420120",
581=> x"8FC5FFF0",
582=> x"20440000",
583=> x"CCA00000",
584=> x"CC800000",
585=> x"D4000177",
586=> x"C8000008",
587=> x"8FC2FFE8",
588=> x"20420001",
589=> x"AFC2FFE8",
590=> x"8FC3FFE8",
591=> x"8FC2000C",
592=> x"00621022",
593=> x"004207D3",
594=> x"10400001",
595=> x"08000235",
596=> x"44800000",
597=> x"048400C0",
598=> x"CC800000",
599=> x"D400017C",
600=> x"C4400000",
601=> x"C8000008",
602=> x"AFC2FFEC",
603=> x"8FC3FFE0",
604=> x"8FC20010",
605=> x"34620000",
606=> x"94600000",
607=> x"8FC20014",
608=> x"00621820",
609=> x"8FC2FFE4",
610=> x"00621020",
611=> x"8FC5FFEC",
612=> x"20440000",
613=> x"CCA00000",
614=> x"CC800000",
615=> x"D4000177",
616=> x"C8000008",
617=> x"8FC2FFE4",
618=> x"20420001",
619=> x"AFC2FFE4",
620=> x"8FC3FFE4",
621=> x"8FC20010",
622=> x"00621022",
623=> x"004207D3",
624=> x"10400001",
625=> x"0800022A",
626=> x"8FC2FFE0",
627=> x"20420001",
628=> x"AFC2FFE0",
629=> x"8FC3FFE0",
630=> x"8FC20008",
631=> x"00621022",
632=> x"004207D3",
633=> x"10400001",
634=> x"08000228",
635=> x"FC000000",
636=> x"D3E00000",
637=> x"C8000038",
638=> x"CC400000",
639=> x"D8000000",
640=> x"C800FFE0",
641=> x"CFE00000",
642=> x"C3C00000",
643=> x"AFC40000",
644=> x"20850000",
645=> x"44800000",
646=> x"048401C8",
647=> x"CCA00000",
648=> x"CC800000",
649=> x"D4000177",
650=> x"C8000008",
651=> x"FC000000",
652=> x"D3E00000",
653=> x"C8000020",
654=> x"CC400000",
655=> x"D8000000",
656=> x"C800FFD8",
657=> x"CFE00000",
658=> x"C3C00000",
659=> x"AFC40000",
660=> x"20820000",
661=> x"8C430000",
662=> x"8FC20000",
663=> x"8C420004",
664=> x"00621025",
665=> x"AFC2FFF0",
666=> x"20450000",
667=> x"44800000",
668=> x"04840180",
669=> x"CCA00000",
670=> x"CC800000",
671=> x"D4000177",
672=> x"C8000008",
673=> x"FC000000",
674=> x"D3E00000",
675=> x"C8000028",
676=> x"CC400000",
677=> x"D8000000",
678=> x"C800FFD8",
679=> x"CFE00000",
680=> x"C3C00000",
681=> x"AFC40000",
682=> x"AFC50004",
683=> x"44800000",
684=> x"04840184",
685=> x"CCA00000",
686=> x"CC800000",
687=> x"D4000177",
688=> x"C8000008",
689=> x"44800000",
690=> x"04840180",
691=> x"CC800000",
692=> x"D400017C",
693=> x"C4400000",
694=> x"C8000008",
695=> x"AFC2FFF0",
696=> x"8FC20000",
697=> x"00430052",
698=> x"8FC2FFF0",
699=> x"00621025",
700=> x"04420400",
701=> x"AFC2FFF4",
702=> x"20450000",
703=> x"44800000",
704=> x"04840180",
705=> x"CCA00000",
706=> x"CC800000",
707=> x"D4000177",
708=> x"C8000008",
709=> x"18000000",
710=> x"FC000000",
711=> x"D3E00000",
712=> x"C8000028",
713=> x"CC400000",
714=> x"D8000000",
715=> x"C800FFD8",
716=> x"CFE00000",
717=> x"C3C00000",
718=> x"AFC40000",
719=> x"20820000",
720=> x"8C430008",
721=> x"8FC20000",
722=> x"8C420004",
723=> x"00621825",
724=> x"8FC20000",
725=> x"8C420000",
726=> x"00621025",
727=> x"AFC2FFF0",
728=> x"20450000",
729=> x"44800000",
730=> x"048401A0",
731=> x"CCA00000",
732=> x"CC800000",
733=> x"D4000177",
734=> x"C8000008",
735=> x"FC000000",
736=> x"D3E00000",
737=> x"C8000028",
738=> x"CC400000",
739=> x"D8000000",
740=> x"C800FFD8",
741=> x"CFE00000",
742=> x"C3C00000",
743=> x"AFC40000",
744=> x"AFC50004",
745=> x"44800000",
746=> x"048401A4",
747=> x"CCA00000",
748=> x"CC800000",
749=> x"D4000177",
750=> x"C8000008",
751=> x"44800000",
752=> x"048401A0",
753=> x"CC800000",
754=> x"D400017C",
755=> x"C4400000",
756=> x"C8000008",
757=> x"AFC2FFF0",
758=> x"04420003",
759=> x"AFC2FFF4",
760=> x"20450000",
761=> x"44800000",
762=> x"048401A0",
763=> x"CCA00000",
764=> x"CC800000",
765=> x"D4000177",
766=> x"C8000008",
767=> x"FC000000",
768=> x"D3E00000",
769=> x"C8000028",
770=> x"CC400000",
771=> x"D8000000",
772=> x"C800FFF8",
773=> x"C3C00000",
774=> x"AFC40000",
775=> x"44600000",
776=> x"04630001",
777=> x"8FC20000",
778=> x"00621016",
779=> x"C8000008",
780=> x"CC400000",
781=> x"D8000000",
782=> x"C0400000",
783=> x"8C430000",
784=> x"8C440004",
785=> x"00640800",
786=> x"CC200000",
787=> x"D8000000",
788=> x"C0400000",
789=> x"8C430000",
790=> x"8C440004",
791=> x"00640802",
792=> x"CC200000",
793=> x"D8000000",
794=> x"C0400000",
795=> x"8C430000",
796=> x"8C440004",
797=> x"00640801",
798=> x"CC200000",
799=> x"D8000000",
800=> x"C0400000",
801=> x"8C430000",
802=> x"8C440004",
803=> x"00640803",
804=> x"CC200000",
805=> x"D8000000",
806=> x"C0400000",
807=> x"8C430000",
808=> x"44808000",
809=> x"00641827",
810=> x"CC600000",
811=> x"D8000000",
812=> x"C800FFE8",
813=> x"C3C00000",
814=> x"AFC40000",
815=> x"20820000",
816=> x"AC0201D8",
817=> x"8C0201DC",
818=> x"AFC2FFF0",
819=> x"C8000018",
820=> x"CC400000",
821=> x"D8000000",
822=> x"C800FFD0",
823=> x"C3C00000",
824=> x"AFC40000",
825=> x"20820000",
826=> x"AFC2FFF0",
827=> x"44400000",
828=> x"04420001",
829=> x"AFC2FFD8",
830=> x"8FC3FFF0",
831=> x"44408000",
832=> x"04420000",
833=> x"00621024",
834=> x"AFC2FFDC",
835=> x"10400001",
836=> x"10000001",
837=> x"08000349",
838=> x"4440FFFF",
839=> x"0442FFFF",
840=> x"AFC2FFD8",
841=> x"8FC2FFF0",
842=> x"004205D8",
843=> x"0C4200FF",
844=> x"AFC2FFE0",
845=> x"2042FF81",
846=> x"AFC2FFE4",
847=> x"8FC2FFF0",
848=> x"20430000",
849=> x"4440007F",
850=> x"04420000",
851=> x"0442FFFF",
852=> x"00621024",
853=> x"AFC2FFE8",
854=> x"20430000",
855=> x"44400080",
856=> x"04420000",
857=> x"00621025",
858=> x"AFC2FFEC",
859=> x"8FC2FFE4",
860=> x"CE000000",
861=> x"0040802A",
862=> x"12000002",
863=> x"D2000000",
864=> x"10000002",
865=> x"D2000000",
866=> x"08000365",
867=> x"20020000",
868=> x"0800037B",
869=> x"8FC2FFE4",
870=> x"54420017",
871=> x"10400001",
872=> x"10000001",
873=> x"08000374",
874=> x"44600000",
875=> x"04630017",
876=> x"8FC2FFE4",
877=> x"00621022",
878=> x"8FC3FFEC",
879=> x"00621817",
880=> x"8FC2FFD8",
881=> x"34620000",
882=> x"94400000",
883=> x"0800037B",
884=> x"8FC2FFE4",
885=> x"2042FFE9",
886=> x"8FC3FFEC",
887=> x"00621816",
888=> x"8FC2FFD8",
889=> x"34620000",
890=> x"94400000",
891=> x"C8000030",
892=> x"CC400000",
893=> x"D8000000",
894=> x"C800FFE0",
895=> x"CFE00000",
896=> x"C3C00000",
897=> x"AFC40000",
898=> x"CC800000",
899=> x"D400038A",
900=> x"C4400000",
901=> x"C8000008",
902=> x"D3E00000",
903=> x"C8000020",
904=> x"CC400000",
905=> x"D8000000",
906=> x"C800FFD8",
907=> x"CFE00000",
908=> x"C3C00000",
909=> x"AFC40000",
910=> x"20820000",
911=> x"CE000000",
912=> x"0040802A",
913=> x"12000002",
914=> x"D2000000",
915=> x"10000002",
916=> x"D2000000",
917=> x"080003A4",
918=> x"8FC20000",
919=> x"00021022",
920=> x"20440000",
921=> x"CC800000",
922=> x"D40003B9",
923=> x"C4400000",
924=> x"C8000008",
925=> x"AFC2FFF0",
926=> x"20430000",
927=> x"44408000",
928=> x"04420000",
929=> x"00621025",
930=> x"AFC2FFF0",
931=> x"080003A9",
932=> x"8FC40000",
933=> x"CC800000",
934=> x"D40003B9",
935=> x"C4400000",
936=> x"C8000008",
937=> x"D3E00000",
938=> x"C8000028",
939=> x"CC400000",
940=> x"D8000000",
941=> x"C800FFE0",
942=> x"CFE00000",
943=> x"C3C00000",
944=> x"AFC40000",
945=> x"CC800000",
946=> x"D40003B9",
947=> x"C4400000",
948=> x"C8000008",
949=> x"D3E00000",
950=> x"C8000020",
951=> x"CC400000",
952=> x"D8000000",
953=> x"C800FFD8",
954=> x"C3C00000",
955=> x"AFC40000",
956=> x"AFC0FFE0",
957=> x"AFC0FFF0",
958=> x"8FC20000",
959=> x"10400001",
960=> x"080003C6",
961=> x"44400000",
962=> x"04420020",
963=> x"AFC2FFEC",
964=> x"8FC2FFF0",
965=> x"08000409",
966=> x"AFC0FFE4",
967=> x"080003D7",
968=> x"8FC30000",
969=> x"8FC2FFE4",
970=> x"00621017",
971=> x"AFC2FFE8",
972=> x"10400001",
973=> x"080003D4",
974=> x"44600000",
975=> x"04630020",
976=> x"8FC2FFE4",
977=> x"00621022",
978=> x"AFC2FFE0",
979=> x"080003DB",
980=> x"8FC2FFE4",
981=> x"20420001",
982=> x"AFC2FFE4",
983=> x"8FC2FFE4",
984=> x"54420020",
985=> x"10400001",
986=> x"080003C8",
987=> x"8FC2FFE0",
988=> x"54420008",
989=> x"10400001",
990=> x"080003F3",
991=> x"8FC2FFE0",
992=> x"2042FFF8",
993=> x"8FC30000",
994=> x"00621016",
995=> x"AFC2FFF0",
996=> x"20430000",
997=> x"4440007F",
998=> x"04420000",
999=> x"0442FFFF",
1000=> x"00621024",
1001=> x"AFC2FFF0",
1002=> x"20430000",
1003=> x"44800000",
1004=> x"0484009E",
1005=> x"8FC2FFE0",
1006=> x"00821022",
1007=> x"004205D2",
1008=> x"00621025",
1009=> x"AFC2FFF0",
1010=> x"08000408",
1011=> x"44600000",
1012=> x"04630008",
1013=> x"8FC2FFE0",
1014=> x"00621022",
1015=> x"8FC30000",
1016=> x"00621017",
1017=> x"AFC2FFF0",
1018=> x"20430000",
1019=> x"4440007F",
1020=> x"04420000",
1021=> x"0442FFFF",
1022=> x"00621024",
1023=> x"AFC2FFF0",
1024=> x"20430000",
1025=> x"44800000",
1026=> x"0484009E",
1027=> x"8FC2FFE0",
1028=> x"00821022",
1029=> x"004205D2",
1030=> x"00621025",
1031=> x"AFC2FFF0",
1032=> x"8FC2FFF0",
1033=> x"C8000028",
1034=> x"CC400000",
1035=> x"D8000000",
1036=> x"C800FFF8",
1037=> x"C3C00000",
1038=> x"AFC40000",
1039=> x"20820000",
1040=> x"AC0201D4",
1041=> x"FC000000",
1042=> x"C8000008",
1043=> x"CC400000",
1044=> x"D8000000",
1045=> x"C800FFE0",
1046=> x"CFE00000",
1047=> x"C3C00000",
1048=> x"44800000",
1049=> x"04840001",
1050=> x"CC800000",
1051=> x"D400040C",
1052=> x"C4400000",
1053=> x"C8000008",
1054=> x"FC000000",
1055=> x"FC000000",
1056=> x"D3E00000",
1057=> x"C8000020",
1058=> x"CC400000",
1059=> x"D8000000",
1060=> x"C800FFE0",
1061=> x"CFE00000",
1062=> x"C3C00000",
1063=> x"44800000",
1064=> x"04840002",
1065=> x"CC800000",
1066=> x"D400040C",
1067=> x"C4400000",
1068=> x"C8000008",
1069=> x"FC000000",
1070=> x"FC000000",
1071=> x"D3E00000",
1072=> x"C8000020",
1073=> x"CC400000",
1074=> x"D8000000",
1075=> x"C800FFE0",
1076=> x"CFE00000",
1077=> x"C3C00000",
1078=> x"AFC40000",
1079=> x"AFC50004",
1080=> x"8FC30000",
1081=> x"8FC20004",
1082=> x"00621025",
1083=> x"04420004",
1084=> x"20440000",
1085=> x"CC800000",
1086=> x"D400040C",
1087=> x"C4400000",
1088=> x"C8000008",
1089=> x"FC000000",
1090=> x"FC000000",
1091=> x"D3E00000",
1092=> x"C8000020",
1093=> x"CC400000",
1094=> x"D8000000",
1095=> x"C800FFE0",
1096=> x"CFE00000",
1097=> x"C3C00000",
1098=> x"AFC40000",
1099=> x"AFC50004",
1100=> x"AFC60008",
1101=> x"8FC30000",
1102=> x"8FC20004",
1103=> x"00621825",
1104=> x"8FC20008",
1105=> x"00621025",
1106=> x"04420008",
1107=> x"20440000",
1108=> x"CC800000",
1109=> x"D400040C",
1110=> x"C4400000",
1111=> x"C8000008",
1112=> x"FC000000",
1113=> x"FC000000",
1114=> x"D3E00000",
1115=> x"C8000020",
1116=> x"CC400000",
1117=> x"D8000000",
1118=> x"C800FFE0",
1119=> x"CFE00000",
1120=> x"C3C00000",
1121=> x"AFC40000",
1122=> x"AFC50004",
1123=> x"8FC30000",
1124=> x"8FC20004",
1125=> x"00621025",
1126=> x"04420010",
1127=> x"20440000",
1128=> x"CC800000",
1129=> x"D400040C",
1130=> x"C4400000",
1131=> x"C8000008",
1132=> x"FC000000",
1133=> x"FC000000",
1134=> x"D3E00000",
1135=> x"C8000020",
1136=> x"CC400000",
1137=> x"D8000000",
1138=> x"C800FFE0",
1139=> x"CFE00000",
1140=> x"C3C00000",
1141=> x"AFC40000",
1142=> x"AFC50004",
1143=> x"AFC60008",
1144=> x"8FC30000",
1145=> x"8FC20004",
1146=> x"00621825",
1147=> x"8FC20008",
1148=> x"00621025",
1149=> x"04420020",
1150=> x"20440000",
1151=> x"CC800000",
1152=> x"D400040C",
1153=> x"C4400000",
1154=> x"C8000008",
1155=> x"FC000000",
1156=> x"FC000000",
1157=> x"D3E00000",
1158=> x"C8000020",
1159=> x"CC400000",
1160=> x"D8000000",
1161=> x"C800FFE0",
1162=> x"CFE00000",
1163=> x"C3C00000",
1164=> x"AFC40000",
1165=> x"20820000",
1166=> x"04420040",
1167=> x"20440000",
1168=> x"CC800000",
1169=> x"D400040C",
1170=> x"C4400000",
1171=> x"C8000008",
1172=> x"FC000000",
1173=> x"FC000000",
1174=> x"D3E00000",
1175=> x"C8000020",
1176=> x"CC400000",
1177=> x"D8000000",
1178=> x"C800FFE0",
1179=> x"CFE00000",
1180=> x"C3C00000",
1181=> x"AFC40000",
1182=> x"20820000",
1183=> x"04420080",
1184=> x"20440000",
1185=> x"CC800000",
1186=> x"D400040C",
1187=> x"C4400000",
1188=> x"C8000008",
1189=> x"FC000000",
1190=> x"FC000000",
1191=> x"D3E00000",
1192=> x"C8000020",
1193=> x"CC400000",
1194=> x"D8000000",
1195=> x"C800FFD8",
1196=> x"CFE00000",
1197=> x"C3C00000",
1198=> x"AFC40000",
1199=> x"AFC50004",
1200=> x"44800000",
1201=> x"04840100",
1202=> x"CC800000",
1203=> x"D400040C",
1204=> x"C4400000",
1205=> x"C8000008",
1206=> x"44800000",
1207=> x"048401D4",
1208=> x"CC800000",
1209=> x"D400017C",
1210=> x"C4400000",
1211=> x"C8000008",
1212=> x"AFC2FFF0",
1213=> x"004201D3",
1214=> x"0C430001",
1215=> x"8FC20000",
1216=> x"AC430000",
1217=> x"8FC2FFF0",
1218=> x"0C43007F",
1219=> x"8FC20004",
1220=> x"AC430000",
1221=> x"FC000000",
1222=> x"FC000000",
1223=> x"D3E00000",
1224=> x"C8000028",
1225=> x"CC400000",
1226=> x"D8000000",
1227=> x"C800FFE0",
1228=> x"CFE00000",
1229=> x"C3C00000",
1230=> x"AFC40000",
1231=> x"20820000",
1232=> x"04420200",
1233=> x"20440000",
1234=> x"CC800000",
1235=> x"D400040C",
1236=> x"C4400000",
1237=> x"C8000008",
1238=> x"FC000000",
1239=> x"FC000000",
1240=> x"D3E00000",
1241=> x"C8000020",
1242=> x"CC400000",
1243=> x"D8000000",
1244=> x"C800FFE0",
1245=> x"CFE00000",
1246=> x"C3C00000",
1247=> x"44800000",
1248=> x"04840300",
1249=> x"CC800000",
1250=> x"D400040C",
1251=> x"C4400000",
1252=> x"C8000008",
1253=> x"44800000",
1254=> x"048401D4",
1255=> x"CC800000",
1256=> x"D400017C",
1257=> x"C4400000",
1258=> x"C8000008",
1259=> x"D3E00000",
1260=> x"C8000020",
1261=> x"CC400000",
1262=> x"D8000000",
1263=> x"C800FFD8",
1264=> x"CFE00000",
1265=> x"C3C00000",
1266=> x"AFC40000",
1267=> x"AFC0FFF0",
1268=> x"080004FE",
1269=> x"8FC2FFF0",
1270=> x"00420092",
1271=> x"8FC30000",
1272=> x"00621020",
1273=> x"8C440000",
1274=> x"CC800000",
1275=> x"D40004CB",
1276=> x"C4400000",
1277=> x"C8000008",
1278=> x"8FC2FFF0",
1279=> x"00420092",
1280=> x"8FC30000",
1281=> x"00621020",
1282=> x"8C420000",
1283=> x"10400001",
1284=> x"080004F5",
1285=> x"FC000000",
1286=> x"D3E00000",
1287=> x"C8000028",
1288=> x"CC400000",
1289=> x"D8000000",
1290=> x"C800FFD8",
1291=> x"CFE00000",
1292=> x"C3C00000",
1293=> x"AFC40000",
1294=> x"44600000",
1295=> x"8C633A58",
1296=> x"44400000",
1297=> x"04420004",
1298=> x"10620001",
1299=> x"08000516",
1300=> x"FC000000",
1301=> x"08000514",
1302=> x"44400000",
1303=> x"8C423A58",
1304=> x"20420001",
1305=> x"44000000",
1306=> x"AC023A58",
1307=> x"00000027",
1308=> x"AFC0FFF0",
1309=> x"0800053D",
1310=> x"44600000",
1311=> x"04630007",
1312=> x"8FC2FFF0",
1313=> x"00621022",
1314=> x"00420092",
1315=> x"8FC30000",
1316=> x"00621017",
1317=> x"0C42000F",
1318=> x"AFC2FFF4",
1319=> x"5442000A",
1320=> x"10400001",
1321=> x"10000001",
1322=> x"08000533",
1323=> x"8FC2FFF4",
1324=> x"20420030",
1325=> x"20440000",
1326=> x"CC800000",
1327=> x"D40004CB",
1328=> x"C4400000",
1329=> x"C8000008",
1330=> x"0800053A",
1331=> x"8FC2FFF4",
1332=> x"20420037",
1333=> x"20440000",
1334=> x"CC800000",
1335=> x"D40004CB",
1336=> x"C4400000",
1337=> x"C8000008",
1338=> x"8FC2FFF0",
1339=> x"20420001",
1340=> x"AFC2FFF0",
1341=> x"8FC2FFF0",
1342=> x"54420008",
1343=> x"10400001",
1344=> x"0800051E",
1345=> x"FC000000",
1346=> x"D3E00000",
1347=> x"C8000028",
1348=> x"CC400000",
1349=> x"D8000000",
1350=> x"C800FF88",
1351=> x"CFE00000",
1352=> x"C3C00000",
1353=> x"AFC40000",
1354=> x"20820000",
1355=> x"AFC2FFDC",
1356=> x"AFC0FFA0",
1357=> x"8FC3FFDC",
1358=> x"44408000",
1359=> x"04420000",
1360=> x"00621024",
1361=> x"AFC2FFC0",
1362=> x"10400001",
1363=> x"10000001",
1364=> x"0800055E",
1365=> x"44800000",
1366=> x"0484002D",
1367=> x"CC800000",
1368=> x"D40004CB",
1369=> x"C4400000",
1370=> x"C8000008",
1371=> x"44400000",
1372=> x"04420001",
1373=> x"AFC2FFA0",
1374=> x"8FC2FFDC",
1375=> x"004205D8",
1376=> x"0C4200FF",
1377=> x"AFC2FFC4",
1378=> x"2042FF81",
1379=> x"0C42FFFF",
1380=> x"AFC2FFC8",
1381=> x"8FC2FFA0",
1382=> x"10400001",
1383=> x"10000001",
1384=> x"0800056E",
1385=> x"8FC3FFDC",
1386=> x"44408000",
1387=> x"04420000",
1388=> x"00621027",
1389=> x"AFC2FFDC",
1390=> x"8FC2FFDC",
1391=> x"AFC2FFA4",
1392=> x"8FC2FFDC",
1393=> x"44A00000",
1394=> x"8CA53A34",
1395=> x"20440000",
1396=> x"CCA00000",
1397=> x"CC800000",
1398=> x"D4000314",
1399=> x"C4400000",
1400=> x"C800000C",
1401=> x"AFC2FFCC",
1402=> x"AFC2FFE0",
1403=> x"CE000000",
1404=> x"0040802A",
1405=> x"12000002",
1406=> x"D2000000",
1407=> x"10000002",
1408=> x"D2000000",
1409=> x"080005A9",
1410=> x"AFC0FFA8",
1411=> x"080005A4",
1412=> x"44A00000",
1413=> x"8CA53A34",
1414=> x"8FC4FFA4",
1415=> x"CCA00000",
1416=> x"CC800000",
1417=> x"D4000314",
1418=> x"C4400000",
1419=> x"C800000C",
1420=> x"AFC2FFD4",
1421=> x"AFC2FFE0",
1422=> x"CE000000",
1423=> x"0040802A",
1424=> x"12000002",
1425=> x"D2000000",
1426=> x"08000598",
1427=> x"D2000000",
1428=> x"8FC2FFA8",
1429=> x"00021022",
1430=> x"AFC2FFA2",
1431=> x"080005E6",
1432=> x"44A00000",
1433=> x"8CA53A50",
1434=> x"8FC4FFA4",
1435=> x"CCA00000",
1436=> x"CC800000",
1437=> x"D400031A",
1438=> x"C4400000",
1439=> x"C800000C",
1440=> x"AFC2FFA4",
1441=> x"8FC2FFA8",
1442=> x"20420001",
1443=> x"AFC2FFA8",
1444=> x"8FC2FFA8",
1445=> x"54420028",
1446=> x"10400001",
1447=> x"08000584",
1448=> x"080005E6",
1449=> x"AFC0FFAC",
1450=> x"080005E2",
1451=> x"44A00000",
1452=> x"8CA53A34",
1453=> x"8FC4FFA4",
1454=> x"CCA00000",
1455=> x"CC800000",
1456=> x"D4000314",
1457=> x"C4400000",
1458=> x"C800000C",
1459=> x"AFC2FFD0",
1460=> x"AFC2FFE0",
1461=> x"8FC2FFAC",
1462=> x"54420028",
1463=> x"10400001",
1464=> x"10000001",
1465=> x"080005D6",
1466=> x"8FC2FFE0",
1467=> x"CE000000",
1468=> x"0040802A",
1469=> x"12000002",
1470=> x"D2000000",
1471=> x"10000002",
1472=> x"D2000000",
1473=> x"080005D6",
1474=> x"8FC3FFE0",
1475=> x"44408000",
1476=> x"04420000",
1477=> x"10620001",
1478=> x"10000001",
1479=> x"080005D6",
1480=> x"44A00000",
1481=> x"8CA53A50",
1482=> x"8FC4FFA4",
1483=> x"CCA00000",
1484=> x"CC800000",
1485=> x"D400031A",
1486=> x"C4400000",
1487=> x"C800000C",
1488=> x"AFC2FFA4",
1489=> x"8FC2FFAC",
1490=> x"2042FFFF",
1491=> x"0C42FFFF",
1492=> x"AFC2FFA2",
1493=> x"080005E6",
1494=> x"44A00000",
1495=> x"8CA53A50",
1496=> x"8FC4FFA4",
1497=> x"CCA00000",
1498=> x"CC800000",
1499=> x"D4000320",
1500=> x"C4400000",
1501=> x"C800000C",
1502=> x"AFC2FFA4",
1503=> x"8FC2FFAC",
1504=> x"20420001",
1505=> x"AFC2FFAC",
1506=> x"8FC2FFAC",
1507=> x"54420028",
1508=> x"10400001",
1509=> x"080005AB",
1510=> x"AFC0FFB0",
1511=> x"08000611",
1512=> x"8FC4FFA4",
1513=> x"CC800000",
1514=> x"D400032C",
1515=> x"C4400000",
1516=> x"C8000008",
1517=> x"20430030",
1518=> x"8FC2FFB0",
1519=> x"00420092",
1520=> x"23C4FFA0",
1521=> x"00821020",
1522=> x"AC430044",
1523=> x"8FC4FFA4",
1524=> x"CC800000",
1525=> x"D400032C",
1526=> x"C4400000",
1527=> x"C8000008",
1528=> x"20440000",
1529=> x"CC800000",
1530=> x"D400037E",
1531=> x"C4400000",
1532=> x"C8000008",
1533=> x"20450000",
1534=> x"8FC4FFA4",
1535=> x"CCA00000",
1536=> x"CC800000",
1537=> x"D4000314",
1538=> x"C4400000",
1539=> x"C800000C",
1540=> x"AFC2FFD8",
1541=> x"44A00000",
1542=> x"8CA53A50",
1543=> x"8FC4FFD8",
1544=> x"CCA00000",
1545=> x"CC800000",
1546=> x"D400031A",
1547=> x"C4400000",
1548=> x"C800000C",
1549=> x"AFC2FFA4",
1550=> x"8FC2FFB0",
1551=> x"20420001",
1552=> x"AFC2FFB0",
1553=> x"8FC2FFB0",
1554=> x"54420002",
1555=> x"10400001",
1556=> x"080005E8",
1557=> x"8FC2FFE4",
1558=> x"04420200",
1559=> x"AC0201D4",
1560=> x"44400000",
1561=> x"0442022E",
1562=> x"AC0201D4",
1563=> x"44400000",
1564=> x"04420001",
1565=> x"AFC2FFB4",
1566=> x"08000629",
1567=> x"8FC2FFB4",
1568=> x"00420092",
1569=> x"23C3FFA0",
1570=> x"00621020",
1571=> x"8C420044",
1572=> x"04420200",
1573=> x"AC0201D4",
1574=> x"8FC2FFB4",
1575=> x"20420001",
1576=> x"AFC2FFB4",
1577=> x"8FC2FFB4",
1578=> x"54420002",
1579=> x"10400001",
1580=> x"0800061F",
1581=> x"44400000",
1582=> x"04420245",
1583=> x"AC0201D4",
1584=> x"8FC2FFA2",
1585=> x"CE000000",
1586=> x"0040802A",
1587=> x"12000002",
1588=> x"D2000000",
1589=> x"10000002",
1590=> x"D2000000",
1591=> x"0800063F",
1592=> x"44400000",
1593=> x"0442022D",
1594=> x"AC0201D4",
1595=> x"8FC2FFA2",
1596=> x"00021022",
1597=> x"0C42FFFF",
1598=> x"AFC2FFA2",
1599=> x"AFC0FFB8",
1600=> x"AFC0FFBC",
1601=> x"0800066E",
1602=> x"8FC3FFA2",
1603=> x"44406666",
1604=> x"04420000",
1605=> x"04426667",
1606=> x"14620000",
1607=> x"B4400000",
1608=> x"00440098",
1609=> x"006207D8",
1610=> x"00822022",
1611=> x"20820000",
1612=> x"00420092",
1613=> x"00441020",
1614=> x"00420052",
1615=> x"00621022",
1616=> x"00430412",
1617=> x"00630418",
1618=> x"8FC2FFBC",
1619=> x"00420092",
1620=> x"23C4FFA0",
1621=> x"00821020",
1622=> x"AC43004C",
1623=> x"8FC2FFA2",
1624=> x"44606666",
1625=> x"04630000",
1626=> x"04636667",
1627=> x"14430000",
1628=> x"B4600000",
1629=> x"00630098",
1630=> x"004207D8",
1631=> x"00621022",
1632=> x"AFC2FFA2",
1633=> x"8FC2FFBC",
1634=> x"00420092",
1635=> x"23C3FFA0",
1636=> x"00621020",
1637=> x"8C42004C",
1638=> x"10400001",
1639=> x"10000001",
1640=> x"0800066B",
1641=> x"8FC2FFBC",
1642=> x"AFC2FFB8",
1643=> x"8FC2FFBC",
1644=> x"20420001",
1645=> x"AFC2FFBC",
1646=> x"8FC2FFBC",
1647=> x"54420002",
1648=> x"10400001",
1649=> x"08000642",
1650=> x"8FC2FFB8",
1651=> x"00420092",
1652=> x"23C3FFA0",
1653=> x"00621020",
1654=> x"8C42004C",
1655=> x"20420030",
1656=> x"04420200",
1657=> x"AC0201D4",
1658=> x"8FC2FFB8",
1659=> x"10400001",
1660=> x"10000001",
1661=> x"08000688",
1662=> x"8FC2FFB8",
1663=> x"2042FFFF",
1664=> x"00420092",
1665=> x"23C3FFA0",
1666=> x"00621020",
1667=> x"8C42004C",
1668=> x"20420030",
1669=> x"04420200",
1670=> x"AC0201D4",
1671=> x"FC000000",
1672=> x"FC000000",
1673=> x"D3E00000",
1674=> x"C8000078",
1675=> x"CC400000",
1676=> x"D8000000",
1677=> x"3F800000",
1678=> x"3ADED289",
1679=> x"C4800000",
1680=> x"3F000000",
1681=> x"461C4000",
1682=> x"40000000",
1683=> x"29E12E13",
1684=> x"41200000",
1685=> x"00000000",
1686=> x"00000000",
1687=> x"00000000",
others=> x"00000000"
	);
	signal rom: memory := initial_value;

	begin
		--output behaviour:
		--necessary turn Auto ROM Replacement on
		process(CLK_A,RST,ADDR_A)
		begin
--			if(RST='1')then
--				ADDR_reg_A <= (others=>'0');
			if(rising_edge(CLK_A))then
--				ADDR_reg_A <= ADDR_A;				
				Q_A <= rom(to_integer(unsigned(ADDR_A)));
			end if;
		end process;
		--surprisingly, the design also works with the synchronous reading logic (ram inferrence)
--		Q_A <= rom(to_integer(unsigned(ADDR_reg_A)));
--		Q_A <= rom(to_integer(unsigned(ADDR_A)));
		
		process(CLK_B,RST,ADDR_B,WREN_B)
		begin
--			if(RST='1')then
--				ADDR_reg_B <= (others=>'0');
--				rom <= initial_value;
--			elsif(rising_edge(CLK) and WREN_B='1')then
			if(rising_edge(CLK_B))then
--				ADDR_reg_B <= ADDR_B;
				if(WREN_B='1')then
					rom(to_integer(unsigned(ADDR_B))) <= D_B;
				end if;
				Q_B <= rom(to_integer(unsigned(ADDR_B)));
			end if;
		end process;		
		--surprisingly, the design also works with the synchronous reading logic (ram inferrence)
--		Q_B <= rom(to_integer(unsigned(ADDR_reg_B)));
--		Q_B <= rom(to_integer(unsigned(ADDR_B)));
end memArch;
